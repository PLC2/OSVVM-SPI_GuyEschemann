package OsvvmTestCommonPkg is
  constant OSVVM_RESULTS_DIR   : string := "" ;
  constant OSVVM_PATH_TO_TESTS : string := "/opt/OsvvmLibraries/" ;
end package OsvvmTestCommonPkg ;
